`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:06:10 04/05/2016 
// Design Name: 
// Module Name:    BlockA 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module BlockA #(parameter nBits=32, parameter M=32, parameter N=16)(
	output [M*N*nBits-1:0]A
    );
assign A={32'h0004b88a,
32'hfffca762,
32'h0005dd12,
32'h00010848,
32'hfffc65e7,
32'h0004342b,
32'hffffcd48,
32'h000612be,
32'h0002afe1,
32'h00049514,
32'hfffb19d0,
32'h00027ebe,
32'h0004dd9b,
32'h00007852,
32'h00018856,
32'h000236da,
32'h0006163e,
32'hfff9314c,
32'h0006e3ae,
32'hffff8a76,
32'h00048043,
32'hfffe5899,
32'hffff09b2,
32'h0007323c,
32'hfffe6ec7,
32'h0001269c,
32'hfffe5d33,
32'h0000963f,
32'h00073d6d,
32'hfffd608f,
32'hfffe4d34,
32'h0002af6d,
32'hfffa67a1,
32'hfff9f4fc,
32'h0000b54f,
32'hfff8adb4,
32'hfffef8a1,
32'hfffc2018,
32'hffff33a6,
32'hffff1543,
32'hfffe02f5,
32'hfffb3e6c,
32'h0004f880,
32'h0002f8ba,
32'h00037428,
32'hfffa159e,
32'h00063d68,
32'h0002096c,
32'h0006335d,
32'h0004da14,
32'hfffa9451,
32'hfffd8e8d,
32'h000628e3,
32'hfffe8f06,
32'hfffd1862,
32'hfffa2ab3,
32'h000751da,
32'hfffc1957,
32'h00048ceb,
32'h00027f78,
32'hfffda87d,
32'h0001aa15,
32'hfff8846c,
32'h0006ad78,
32'h0001fc42,
32'h0002ec24,
32'hfffabd4a,
32'hfffaeec8,
32'hfffb3a4b,
32'hfff9f263,
32'h000020ac,
32'hfffc5ef8,
32'hfff910eb,
32'h0005cc35,
32'hfff96836,
32'hfffb2c07,
32'h000142d4,
32'h00042e9a,
32'hffff6fce,
32'hfffba24f,
32'hfff9f68e,
32'hfffd41a9,
32'hfffc5cd5,
32'h00046a0d,
32'hfffc7501,
32'hfffa7ac7,
32'h0000295d,
32'hfffea17c,
32'h0005c70c,
32'hfff8ee1c,
32'hfffe7d26,
32'hfffa6b93,
32'hfffa1dd5,
32'hfffeda0f,
32'hfffedd80,
32'h000323a4,
32'hfffcad6f,
32'h0006c0da,
32'h00051c5b,
32'hfffd2b11,
32'hfffaaedf,
32'h0006a179,
32'h0004c3b1,
32'h00016c67,
32'h00063305,
32'hffffd939,
32'h00006734,
32'h00077c78,
32'h00061839,
32'hfff9dcc3,
32'hffff69eb,
32'hfffc0b20,
32'h0000b406,
32'hfff90446,
32'hfffc5072,
32'h00006d91,
32'hfffa8a81,
32'h0006d78e,
32'h00046c27,
32'hfffc6ee5,
32'h00047159,
32'hfffb04d7,
32'hfffec083,
32'hfffb111b,
32'h0005b1df,
32'hfffc7f40,
32'h00040d6a,
32'hfffa4a7b,
32'h0006dcd4,
32'hffff14c7,
32'h0004b6db,
32'hfffafc17,
32'h00058a15,
32'h000120cd,
32'h00022a2e,
32'h00018aeb,
32'hfff9fb0e,
32'h00072e22,
32'h00025a58,
32'hfff8fd30,
32'h0004c433,
32'hffface0b,
32'hfffd564b,
32'h00019c0c,
32'h0006f92c,
32'hfffe392f,
32'hfffc2723,
32'h0001879c,
32'h00013211,
32'hfff9658e,
32'hfffe2ddc,
32'h00032b12,
32'hfffc6d96,
32'h000330bf,
32'h0001eb6b,
32'h0000eb02,
32'hfffc6932,
32'hfffcb70f,
32'h00044566,
32'hffff4087,
32'hfffadd3c,
32'h0003fb96,
32'h0006705f,
32'hfffc71cf,
32'h0000bf77,
32'hfffc058e,
32'h0004ac78,
32'hfffbd382,
32'hfffd87c5,
32'h000001d0,
32'hfffce138,
32'h0005ba5e,
32'h00016a54,
32'hffff19ed,
32'hffff9203,
32'hffff6182,
32'h00070f14,
32'h00046d91,
32'hfffdbff0,
32'h00024faa,
32'hfffaaca0,
32'hfffdcc21,
32'h00007e0d,
32'hfffa42e2,
32'h0002b228,
32'hffff90fb,
32'hfffef98a,
32'h000289a2,
32'hfff8d673,
32'h0000683a,
32'hfff90954,
32'h00026dde,
32'h0006db85,
32'hfffb4d97,
32'hfffb72ed,
32'h0002d695,
32'h00054ba4,
32'h0004d163,
32'hfffdc2cb,
32'hfffcf33c,
32'hfffa8c5d,
32'hfff964f0,
32'hfff8bb78,
32'hfffb5b44,
32'hfffee0ff,
32'hffff5c82,
32'hfffb235c,
32'h00040de5,
32'hffffc7d8,
32'hffffd8b2,
32'hfffc4429,
32'h0003b8e7,
32'h0001d4b1,
32'hfff8bb26,
32'h000695c4,
32'hfffd481c,
32'h00035183,
32'h0002bac6,
32'h000742ce,
32'hfffe08a4,
32'hfffd30d7,
32'h0005a16d,
32'h0003538d,
32'hfffdc0d6,
32'h00048114,
32'hffff2f0d,
32'h0001bd9d,
32'hffff4214,
32'hfffdc3a8,
32'hfff92536,
32'h0005a39f,
32'hfffedccd,
32'hfffa19f7,
32'hfff922f0,
32'hfffb01ed,
32'hffff6930,
32'hfffaec1a,
32'h00004552,
32'hffff9a30,
32'h00026e1e,
32'hfffaa0d8,
32'h000231d8,
32'hffff996e,
32'hfff9c1e0,
32'h000032e1,
32'hfffb08ec,
32'h0000c09a,
32'h00001e2d,
32'h00024e6e,
32'hfff9925a,
32'hfffa17df,
32'h0007397d,
32'hfffb2e76,
32'h0006a783,
32'hfffaca73,
32'hfffebe0d,
32'hfffed390,
32'h000323f6,
32'hfffdc65f,
32'hfffbef46,
32'hfffe86f1,
32'h00023c9a,
32'h0001d64e,
32'hfff9c861,
32'hffffe9a1,
32'h00005323,
32'hfffe160e,
32'hfffad898,
32'hfffed7e2,
32'h000210ce,
32'hfffd9deb,
32'h00052102,
32'h00063c6d,
32'h0003d1ff,
32'h0004f662,
32'h00063337,
32'hfff9a3b6,
32'h000379d0,
32'h00014e40,
32'hfffc6fef,
32'h00042f8f,
32'hfff9f371,
32'hfffb78c6,
32'h00055535,
32'hfff9e9d7,
32'h0006dd8b,
32'h00019c60,
32'h0004fe67,
32'h00046213,
32'hfffca3f0,
32'h0001476a,
32'hfffac922,
32'hfffc1947,
32'h00023758,
32'hfffb9dbb,
32'h000483e5,
32'h000339be,
32'h0004c5b1,
32'hffffd867,
32'h00022be5,
32'h00017a55,
32'hfffc1c51,
32'hfffb604d,
32'hfffc58bc,
32'h0006e473,
32'h0002b20f,
32'h0000bef0,
32'h0004e323,
32'hfffa598b,
32'hffff438c,
32'hfffd04c9,
32'hfff8f035,
32'h00060e49,
32'h0004c361,
32'hfffd97a8,
32'hfffe24e3,
32'hffff9059,
32'h0002a44f,
32'h0003938f,
32'h0001b3b0,
32'h0002560b,
32'h00025394,
32'h00064206,
32'h0000933c,
32'hfffb4235,
32'h0000b484,
32'hffff9058,
32'h00066ecd,
32'h0005dd24,
32'h0003562b,
32'h0006c643,
32'hfffb5d26,
32'h0002f072,
32'hfffcd602,
32'hfffc248b,
32'h00013bd6,
32'hfff90922,
32'hfffaf06e,
32'hfffcc99f,
32'h00077128,
32'hfffc196b,
32'hfffcf1df,
32'hfffbf513,
32'h00037478,
32'hfffd8330,
32'hfffabf7c,
32'h00064e13,
32'hfffeec7e,
32'h0002ff92,
32'h000293be,
32'h000642e9,
32'h00009c70,
32'h00053ca8,
32'hfffa48f3,
32'h0003dba6,
32'hfff9ac32,
32'hfffec24e,
32'h0003ab9f,
32'h00052a25,
32'hffffd442,
32'h0002fb2f,
32'h000264e2,
32'hfff94a48,
32'hffffbaf7,
32'h000213f5,
32'h0002ed57,
32'hfffc8932,
32'h00058c93,
32'h00068289,
32'hfffff9b8,
32'h0003ce52,
32'hffff23e2,
32'hfff93eac,
32'hfffb5596,
32'hfffb6be5,
32'h00012d89,
32'hfffb7797,
32'h00004768,
32'h00039160,
32'hfffa4f26,
32'hfff9010a,
32'hfff98518,
32'h0003fb85,
32'hfffc78c0,
32'h0002ae58,
32'h0006e56b,
32'hfffe34e9,
32'hfffa198c,
32'h00060a6e,
32'h0002cd38,
32'hfffbe38a,
32'hfffc0f2b,
32'hfff8f547,
32'h00071839,
32'hfffc896b,
32'h000157b5,
32'hfff98837,
32'hfffc5265,
32'hfffb5476,
32'hfffd4568,
32'h0003ddb9,
32'hfffd9b15,
32'h0001046f,
32'h0006edb0,
32'h0006abfc,
32'hfffb40af,
32'hfffb0f85,
32'hffff61fb,
32'h0003a93f,
32'h00023c21,
32'hfffed7b0,
32'hfffbe490,
32'hfffd4b43,
32'hfffbdc50,
32'hfffccffe,
32'hfffa49c9,
32'h0003a5a1,
32'h0001476e,
32'hfff9a348,
32'hfff891cc,
32'hffffdceb,
32'hfffe06fb,
32'hfffbea3b,
32'h0006f243,
32'h00000016,
32'h00048145,
32'h0000b7d3,
32'hfffe44f0,
32'h00007685,
32'h0002847a,
32'hfff9dde0,
32'h000698f2,
32'hfffe6227,
32'hfffbdb70,
32'hfff94f2b,
32'h00041fa8,
32'hffffd6bb,
32'h0001e260,
32'hffff0915,
32'h0000b3bc,
32'hffffb2e7,
32'hffff4e95,
32'h0006a41c,
32'h00013eab,
32'h00025112,
32'h00052a77,
32'h000124a5,
32'h00022eeb,
32'h00025509,
32'h0003c4de,
32'h00007643,
32'h0004c272,
32'hfffd90d8,
32'h00043413,
32'hfffd2aa2,
32'h00005129,
32'h00061222,
32'hfffefc62,
32'hfffec423,
32'hfffc46ef,
32'hfffe9d42,
32'hfffdaabc,
32'h0002c01d,
32'hffffb124,
32'hfffb115b,
32'hfffc5391,
32'h00043001,
32'h000587ca,
32'h00060035,
32'hfff9b786,
32'h000659c7,
32'hfffbf953,
32'h0001a5e3,
32'h0004e134,
32'h00073eec,
32'hfffcdb4b,
32'h0004ccba,
32'h00043532,
32'h0000b2eb,
32'h000216fa,
32'h00031738,
32'h000016e0,
32'h0006829a,
32'hfff9c43c,
32'hfffe09e8,
32'h000670d8,
32'hfffef3ff,
32'hffffd55e,
32'h0001c3d7,
32'hfff9c086,
32'hfffd0596,
32'h0001c1a1,
32'h00034680,
32'h0002a146,
32'hfffee2cc,
32'h0000abb6,
32'hfff8fa3d,
32'h0002fc74,
32'hfffa72d7,
32'hfffe7f2a,
32'hfffa2b05,
32'h000422bd,
32'hfffb45b2,
32'h0001dc64,
32'h00056442,
32'hfffa7f60,
32'h00030438,
32'hfffc7aae,
32'h0007079d,
32'hfff899c9,
32'h00022aa9,
32'h000235ad
};
endmodule
